netcdf mesonet {
dimensions:
	recNum = UNLIMITED ;
	maxStaTypeLen = 11 ;
	maxStaIdLen = 6 ;
	maxNameLength = 51 ;
	maxSensor = 2 ;
	QCcheckNum = 10 ;
	dateTimeLen = 23 ;
variables:
	char stationId(recNum, maxStaIdLen) ;
		stationId:long_name = "alphanumeric station Id" ;
		stationId:reference = "station table" ;
	char stationType(recNum, maxStaTypeLen) ;
		stationType:long_name = "LDAD station type" ;
	char stationName(recNum, maxNameLength) ;
		stationName:long_name = "alphanumeric station name" ;
		stationName:reference = "station table" ;
	float latitude(recNum) ;
		latitude:long_name = "latitude" ;
		latitude:units = "degree_north" ;
		latitude:_FillValue = 3.402823e+38f ;
		latitude:missing_value = -9999.f ;
		latitude:reference = "station table" ;
		latitude:standard_name = "latitude" ;
	float longitude(recNum) ;
		longitude:long_name = "longitude" ;
		longitude:units = "degree_east" ;
		longitude:_FillValue = 3.402823e+38f ;
		longitude:missing_value = -9999.f ;
		longitude:reference = "station table" ;
		longitude:standard_name = "longitude" ;
	float elevation(recNum) ;
		elevation:long_name = "elevation" ;
		elevation:units = "meter" ;
		elevation:_FillValue = 3.402823e+38f ;
		elevation:missing_value = -9999.f ;
		elevation:reference = "station table" ;
		elevation:standard_name = "elevation" ;
	double observationTime(recNum) ;
		observationTime:long_name = "time of observation" ;
		observationTime:units = "seconds since 1970-1-1 00:00:00.0" ;
		observationTime:_FillValue = 3.40282346e+38 ;
		observationTime:missing_value = -9999. ;
		observationTime:standard_name = "time" ;
	float stationPressure(recNum) ;
		stationPressure:long_name = "station pressure" ;
		stationPressure:units = "pascal" ;
		stationPressure:_FillValue = 3.402823e+38f ;
		stationPressure:missing_value = -9999.f ;
		stationPressure:standard_name = "surface_air_pressure" ;
	float temperature(recNum) ;
		temperature:long_name = "temperature" ;
		temperature:units = "kelvin" ;
		temperature:_FillValue = 3.402823e+38f ;
		temperature:missing_value = -9999.f ;
		temperature:standard_name = "air_temperature" ;
	int temperatureQCR(recNum) ;
		temperatureQCR:long_name = "Temperature QC Results word" ;
		temperatureQCR:NoBitsSet = "No QC failures" ;
		temperatureQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		temperatureQCR:Bit2Set = "Validity check failed" ;
		temperatureQCR:Bit3Set = "Reserved" ;
		temperatureQCR:Bit4Set = "Internal Consistency check failed" ;
		temperatureQCR:Bit5Set = "Temporal Consistency check failed" ;
		temperatureQCR:Bit6Set = "Statistical Spatial Consistency check failed" ;
		temperatureQCR:Bit7Set = "Spatial Consistency check failed" ;
		temperatureQCR:Bit8Set = "Forecast Model Consistency check failed" ;
		temperatureQCR:Bit9Set = "Reserved" ;
		temperatureQCR:Bit10Set = "Kalman Filter failed" ;
		temperatureQCR:reference = "Global Attributes Section" ;
	float temperatureQCD(recNum, QCcheckNum) ;
		temperatureQCD:long_name = "temperature QC departures" ;
		temperatureQCD:_FillValue = 3.402823e+38f ;
		temperatureQCD:units = "kelvin" ;
		temperatureQCD:pos1 = "Average ob departure from QC check estimates" ;
		temperatureQCD:pos2 = "Reserved" ;
		temperatureQCD:pos3 = "Reserved" ;
		temperatureQCD:pos4 = "Internal consistency check departure" ;
		temperatureQCD:pos5 = "Temporal consistency departure" ;
		temperatureQCD:pos6 = "Reserved" ;
		temperatureQCD:pos7 = "Spatial consistency departure" ;
		temperatureQCD:pos8 = "Model consistency departure" ;
		temperatureQCD:pos9 = "Reserved" ;
		temperatureQCD:pos10 = "Kalman filter departure" ;
		temperatureQCD:reference = "Global Attributes Section" ;
	float dewpoint(recNum) ;
		dewpoint:long_name = "dew point temperature" ;
		dewpoint:units = "kelvin" ;
		dewpoint:_FillValue = 3.402823e+38f ;
		dewpoint:missing_value = -9999.f ;
		dewpoint:standard_name = "dew_point_temperature" ;
	int dewpointQCR(recNum) ;
		dewpointQCR:long_name = "dew point QC results word" ;
		dewpointQCR:NoBitsSet = "No QC failures" ;
		dewpointQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		dewpointQCR:Bit2Set = "Validity check failed" ;
		dewpointQCR:Bit3Set = "Reserved" ;
		dewpointQCR:Bit4Set = "Internal Consistency check failed" ;
		dewpointQCR:Bit5Set = "Temporal Consistency check failed" ;
		dewpointQCR:Bit6Set = "Statistical Spatial Consistency check failed" ;
		dewpointQCR:Bit7Set = "Spatial Consistency check failed" ;
		dewpointQCR:Bit8Set = "Forecast Model Consistency check failed" ;
		dewpointQCR:reference = "Global Attributes Section" ;
	float dewpointQCD(recNum, QCcheckNum) ;
		dewpointQCD:long_name = "dew point QC departures" ;
		dewpointQCD:_FillValue = 3.402823e+38f ;
		dewpointQCD:units = "kelvin" ;
		dewpointQCD:pos1 = "Average ob departure from QC check estimates" ;
		dewpointQCD:pos2 = "Reserved" ;
		dewpointQCD:pos3 = "Reserved" ;
		dewpointQCD:pos4 = "Internal consistency check departure" ;
		dewpointQCD:pos5 = "Temporal consistency check departure" ;
		dewpointQCD:pos6 = "Reserved" ;
		dewpointQCD:pos7 = "Spatial consistency check departure" ;
		dewpointQCD:pos8 = "Forecast Model consistency check departure" ;
		dewpointQCD:reference = "Global Attributes Section" ;
	float relHumidity(recNum) ;
		relHumidity:long_name = "relative humidity" ;
		relHumidity:units = "percent" ;
		relHumidity:_FillValue = 3.402823e+38f ;
		relHumidity:missing_value = -9999.f ;
		relHumidity:standard_name = "relative_humidity" ;
	float windDir(recNum) ;
		windDir:long_name = "wind direction" ;
		windDir:units = "degree" ;
		windDir:_FillValue = 3.402823e+38f ;
		windDir:missing_value = -9999.f ;
		windDir:standard_name = "wind_from_direction" ;
	int windDirQCR(recNum) ;
		windDirQCR:long_name = "wind direction QC results word" ;
		windDirQCR:NoBitsSet = "No QC failures" ;
		windDirQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		windDirQCR:Bit2Set = "Validity check failed" ;
		windDirQCR:Bit3Set = "Reserved" ;
		windDirQCR:Bit4Set = "Internal Consistency check failed" ;
		windDirQCR:Bit5Set = "Temporal Consistency check failed" ;
		windDirQCR:Bit6Set = "Statistical Spatial Consistency check failed" ;
		windDirQCR:Bit7Set = "Spatial Consistency check failed" ;
		windDirQCR:Bit8Set = "Forecast Model Consistency check failed" ;
		windDirQCR:reference = "Global Attributes Section" ;
	float windDirQCD(recNum, QCcheckNum) ;
		windDirQCD:long_name = "wind direction QC departures" ;
		windDirQCD:units = "degree" ;
		windDirQCD:_FillValue = 3.402823e+38f ;
		windDirQCD:pos1 = "Average ob departure from QC check estimates" ;
		windDirQCD:pos2 = "Reserved" ;
		windDirQCD:pos3 = "Reserved" ;
		windDirQCD:pos4 = "Internal Consistency check departure" ;
		windDirQCD:pos5 = "Temporal Consistency check departure" ;
		windDirQCD:pos6 = "Reserved" ;
		windDirQCD:pos7 = "Spatial Consistency check departure" ;
		windDirQCD:pos8 = "Forecast Model Consistency check departure" ;
		windDirQCD:reference = "Global Attributes Section" ;
	float windSpeed(recNum) ;
		windSpeed:long_name = "wind speed" ;
		windSpeed:units = "meter/sec" ;
		windSpeed:_FillValue = 3.402823e+38f ;
		windSpeed:missing_value = -9999.f ;
		windSpeed:valid_min = 0. ;
		windSpeed:standard_name = "wind_speed" ;
	int windSpeedQCR(recNum) ;
		windSpeedQCR:long_name = "wind speed QC results word" ;
		windSpeedQCR:NoBitsSet = "No QC failures" ;
		windSpeedQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		windSpeedQCR:Bit2Set = "Validity check failed" ;
		windSpeedQCR:Bit3Set = "Reserved" ;
		windSpeedQCR:Bit4Set = "Internal Consistency check failed" ;
		windSpeedQCR:Bit5Set = "Temporal Consistency check failed" ;
		windSpeedQCR:Bit6Set = "Statistical Spatial Consistency check failed" ;
		windSpeedQCR:Bit7Set = "Spatial Consistency check failed" ;
		windSpeedQCR:Bit8Set = "Forecast Model Consistency check failed" ;
		windSpeedQCR:reference = "Global Attributes Section" ;
	float windSpeedQCD(recNum, QCcheckNum) ;
		windSpeedQCD:long_name = "wind speed QC departures" ;
		windSpeedQCD:units = "meter/sec" ;
		windSpeedQCD:_FillValue = 3.402823e+38f ;
		windSpeedQCD:pos1 = "Average ob departure from QC check estimates" ;
		windSpeedQCD:pos2 = "Reserved" ;
		windSpeedQCD:pos3 = "Reserved" ;
		windSpeedQCD:pos4 = "Internal Consistency check departure" ;
		windSpeedQCD:pos5 = "Temporal Consistency check departure" ;
		windSpeedQCD:pos6 = "Reserved" ;
		windSpeedQCD:pos7 = "Spatial Consistency check departure" ;
		windSpeedQCD:pos8 = "Forecast Model Consistency check departure" ;
		windSpeedQCD:reference = "Global Attributes Section" ;
	float windGust(recNum) ;
		windGust:long_name = "wind gust" ;
		windGust:units = "meter/sec" ;
		windGust:_FillValue = 3.402823e+38f ;
		windGust:missing_value = -9999.f ;
		windGust:valid_min = 0. ;
		windGust:standard_name = "wind_gust" ;
	float windDirMax(recNum) ;
		windDirMax:long_name = "wind direction at gust" ;
		windDirMax:units = "degree" ;
		windDirMax:_FillValue = 3.402823e+38f ;
		windDirMax:missing_value = -9999.f ;
		windDirMax:standard_name = "wind_gust_from_direction" ;
	float visibility(recNum) ;
		visibility:long_name = "visibility" ;
		visibility:units = "meter" ;
		visibility:_FillValue = 3.402823e+38f ;
		visibility:missing_value = -9999.f ;
		visibility:valid_min = 0. ;
		visibility:standard_name = "visibility_in_air" ;
	int visibilityQCR(recNum) ;
		visibilityQCR:long_name = "visibility QC results word" ;
		visibilityQCR:NoBitsSet = "No QC failures" ;
		visibilityQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		visibilityQCR:Bit2Set = "Validity check failed" ;
		visibilityQCR:Bit3Set = "Reserved" ;
		visibilityQCR:Bit4Set = "Internal Consistency check failed" ;
		visibilityQCR:Bit5Set = "Reserved" ;
		visibilityQCR:Bit6Set = "Statistical Spatial Consistency check failed" ;
		visibilityQCR:Bit7Set = "Spatial Consistency check failed" ;
		visibilityQCR:Bit8Set = "Forecast Model Consistency check failed" ;
		visibilityQCR:reference = "Global Attributes Section" ;
	float visibilityQCD(recNum, QCcheckNum) ;
		visibilityQCD:long_name = "visibility QC departures" ;
		visibilityQCD:units = "meter" ;
		visibilityQCD:_FillValue = 3.402823e+38f ;
		visibilityQCD:pos1 = "Average ob departure from QC check estimates" ;
		visibilityQCD:pos2 = "Reserved" ;
		visibilityQCD:pos3 = "Reserved" ;
		visibilityQCD:pos4 = "Internal Consistency check departure" ;
		visibilityQCD:pos5 = "Reserved" ;
		visibilityQCD:pos6 = "Reserved" ;
		visibilityQCD:pos7 = "Spatial Consistency check departure" ;
		visibilityQCD:pos8 = "Forecast Model Consistency check departure" ;
		visibilityQCD:reference = "Global Attributes Section" ;
	float precipAccum(recNum) ;
		precipAccum:long_name = "precip accumulation" ;
		precipAccum:units = "mm" ;
		precipAccum:_FillValue = 3.402823e+38f ;
		precipAccum:missing_value = -9999.f ;
	int precipAccumQCR(recNum) ;
		precipAccumQCR:long_name = "precip amount QC results word" ;
		precipAccumQCR:NoBitsSet = "No QC failures" ;
		precipAccumQCR:Bit1Set = "Master-at least 1 check failed" ;
		precipAccumQCR:Bit2Set = "Validity check failed" ;
		precipAccumQCR:Bit3Set = "Reserved" ;
		precipAccumQCR:Bit4Set = "Internal Consistency check failed" ;
		precipAccumQCR:reference = "Global Attributes Section" ;
	float precipAccumQCD(recNum, QCcheckNum) ;
		precipAccumQCD:long_name = "precip amount QC departures" ;
		precipAccumQCD:units = "mm" ;
		precipAccumQCD:_FillValue = 3.402823e+38f ;
		precipAccumQCD:pos1 = "Average ob departure" ;
		precipAccumQCD:pos2 = "Reserved" ;
		precipAccumQCD:pos3 = "Reserved" ;
		precipAccumQCD:pos4 = "Internal Consistency check departure" ;
		precipAccumQCD:reference = "Global Attributes Section" ;
	float precipRate(recNum) ;
		precipRate:long_name = "precipitation rate" ;
		precipRate:units = "meter/second" ;
		precipRate:_FillValue = 3.402823e+38f ;
		precipRate:missing_value = -9999.f ;
		precipRate:standard_name = "rainfall_rate" ;
	short precipType(recNum, maxSensor) ;
		precipType:long_name = "precipitation type" ;
		precipType:value0 = "no precipitation" ;
		precipType:value1 = "precipitation present but unclassified" ;
		precipType:value2 = "rain" ;
		precipType:value3 = "snow" ;
		precipType:value4 = "mixed rain and snow" ;
		precipType:value5 = "light" ;
		precipType:value6 = "light freezing" ;
		precipType:value7 = "freezing rain" ;
		precipType:value8 = "sleet" ;
		precipType:value9 = "hail" ;
		precipType:value10 = "other" ;
		precipType:value11 = "unidentified" ;
		precipType:value12 = "unknown" ;
		precipType:value13 = "frozen" ;
		precipType:value14 = "ice pellets" ;
		precipType:value15 = "recent" ;
		precipType:value16 = "lens dirty" ;
		precipType:value29 = "RPU-to-maxSensor communications failure" ;
		precipType:value30 = "sensor failure" ;
		precipType:_FillValue = -32767s ;
		precipType:missing_value = -9999s ;
	short precipIntensity(recNum, maxSensor) ;
		precipIntensity:long_name = "precipitation intensity" ;
		precipIntensity:value0 = "precipitation intensity info not available" ;
		precipIntensity:value1 = "none" ;
		precipIntensity:value2 = "light" ;
		precipIntensity:value3 = "moderate" ;
		precipIntensity:value4 = "heavy" ;
		precipIntensity:value5 = "slight" ;
		precipIntensity:value6 = "other" ;
		precipIntensity:_FillValue = -32767s ;
		precipIntensity:missing_value = -9999s ;
	double timeSinceLastPcp(recNum) ;
		timeSinceLastPcp:long_name = "time since last precip" ;
		timeSinceLastPcp:units = "second" ;
		timeSinceLastPcp:_FillValue = 3.40282346e+38 ;
		timeSinceLastPcp:valid_min = 0 ;
		timeSinceLastPcp:missing_value = -9999. ;
	float solarRadiation(recNum) ;
		solarRadiation:long_name = "solar radiation" ;
		solarRadiation:units = "watt/meter2" ;
		solarRadiation:_FillValue = 3.402823e+38f ;
		solarRadiation:missing_value = -9999.f ;
	float roadSurfaceFriction1(recNum) ;
		roadSurfaceFriction1:long_name = "Road surface friction" ;
		roadSurfaceFriction1:units = "percent" ;
		roadSurfaceFriction1:_FillValue = 3.402823e+38f ;
		roadSurfaceFriction1:missing_value = -9999.f ;
	short roadState1(recNum) ;
		roadState1:long_name = "Road State - sensor 1" ;
		roadState1:value0 = "No report" ;
		roadState1:value1 = "Dry" ;
		roadState1:value2 = "Moist" ;
		roadState1:value3 = "Moist and chemically treated" ;
		roadState1:value4 = "Wet" ;
		roadState1:value5 = "Wet and chemically treated" ;
		roadState1:value6 = "Ice" ;
		roadState1:value7 = "Frost" ;
		roadState1:value8 = "Snow" ;
		roadState1:value9 = "Snow/Ice Watch" ;
		roadState1:value10 = "Snow/Ice Warning" ;
		roadState1:value11 = "Wet Above Freezing" ;
		roadState1:value12 = "Wet Below Freezing" ;
		roadState1:value13 = "Absorption" ;
		roadState1:value14 = "Absorption at Dewpoint" ;
		roadState1:value15 = "Dew" ;
		roadState1:value16 = "Black Ice Warning" ;
		roadState1:value17 = "Other" ;
		roadState1:value18 = "Slush" ;
		roadState1:_FillValue = -32767s ;
		roadState1:missing_value = -9999 ;
	short roadState2(recNum) ;
		roadState2:long_name = "Road State - sensor 2" ;
		roadState2:value0 = "No report" ;
		roadState2:value1 = "Dry" ;
		roadState2:value2 = "Moist" ;
		roadState2:value3 = "Moist and chemically treated" ;
		roadState2:value4 = "Wet" ;
		roadState2:value5 = "Wet and chemically treated" ;
		roadState2:value6 = "Ice" ;
		roadState2:value7 = "Frost" ;
		roadState2:value8 = "Snow" ;
		roadState2:value9 = "Snow/Ice Watch" ;
		roadState2:value10 = "Snow/Ice Warning" ;
		roadState2:value11 = "Wet Above Freezing" ;
		roadState2:value12 = "Wet Below Freezing" ;
		roadState2:value13 = "Absorption" ;
		roadState2:value14 = "Absorption at Dewpoint" ;
		roadState2:value15 = "Dew" ;
		roadState2:value16 = "Black Ice Warning" ;
		roadState2:value17 = "Other" ;
		roadState2:value18 = "Slush" ;
		roadState2:_FillValue = -32767s ;
		roadState2:missing_value = -9999 ;
	short roadState3(recNum) ;
		roadState3:long_name = "Road State - sensor 3" ;
		roadState3:value0 = "No report" ;
		roadState3:value1 = "Dry" ;
		roadState3:value2 = "Moist" ;
		roadState3:value3 = "Moist and chemically treated" ;
		roadState3:value4 = "Wet" ;
		roadState3:value5 = "Wet and chemically treated" ;
		roadState3:value6 = "Ice" ;
		roadState3:value7 = "Frost" ;
		roadState3:value8 = "Snow" ;
		roadState3:value9 = "Snow/Ice Watch" ;
		roadState3:value10 = "Snow/Ice Warning" ;
		roadState3:value11 = "Wet Above Freezing" ;
		roadState3:value12 = "Wet Below Freezing" ;
		roadState3:value13 = "Absorption" ;
		roadState3:value14 = "Absorption at Dewpoint" ;
		roadState3:value15 = "Dew" ;
		roadState3:value16 = "Black Ice Warning" ;
		roadState3:value17 = "Other" ;
		roadState3:value18 = "Slush" ;
		roadState3:_FillValue = -32767s ;
		roadState3:missing_value = -9999 ;
	float roadTemperature1(recNum) ;
		roadTemperature1:long_name = "Road temperature - sensor 1" ;
		roadTemperature1:units = "kelvin" ;
		roadTemperature1:_FillValue = 3.402823e+38f ;
		roadTemperature1:missing_value = -9999.f ;
		roadTemperature1:standard_name = "pavement_temperature" ;
	float roadTemperature2(recNum) ;
		roadTemperature2:long_name = "Road temperature - sensor 2" ;
		roadTemperature2:units = "kelvin" ;
		roadTemperature2:_FillValue = 3.402823e+38f ;
		roadTemperature2:missing_value = -9999.f ;
	float roadTemperature3(recNum) ;
		roadTemperature3:long_name = "Road temperature - sensor 3" ;
		roadTemperature3:units = "kelvin" ;
		roadTemperature3:_FillValue = 3.402823e+38f ;
		roadTemperature3:missing_value = -9999.f ;
	float roadTemperature4(recNum) ;
		roadTemperature4:long_name = "Road temperature - sensor 4" ;
		roadTemperature4:units = "kelvin" ;
		roadTemperature4:_FillValue = 3.402823e+38f ;
		roadTemperature4:missing_value = -9999.f ;
	float roadSubsurfaceTemp1(recNum) ;
		roadSubsurfaceTemp1:long_name = "Road subsurface temp - sensor 1" ;
		roadSubsurfaceTemp1:units = "kelvin" ;
		roadSubsurfaceTemp1:_FillValue = 3.402823e+38f ;
		roadSubsurfaceTemp1:missing_value = -9999.f ;
	float roadSubsurfaceTemp2(recNum) ;
		roadSubsurfaceTemp2:long_name = "Road subsurface temp - sensor 2" ;
		roadSubsurfaceTemp2:units = "kelvin" ;
		roadSubsurfaceTemp2:_FillValue = 3.402823e+38f ;
		roadSubsurfaceTemp2:missing_value = -9999.f ;
	float roadSubsurfaceTemp3(recNum) ;
		roadSubsurfaceTemp3:long_name = "Road subsurface temp - sensor 3" ;
		roadSubsurfaceTemp3:units = "kelvin" ;
		roadSubsurfaceTemp3:_FillValue = 3.402823e+38f ;
		roadSubsurfaceTemp3:missing_value = -9999.f ;
	float roadSubsurfaceTemp4(recNum) ;
		roadSubsurfaceTemp4:long_name = "Road subsurface temp - sensor 4" ;
		roadSubsurfaceTemp4:units = "kelvin" ;
		roadSubsurfaceTemp4:_FillValue = 3.402823e+38f ;
		roadSubsurfaceTemp4:missing_value = -9999.f ;
	float roadIceDepth1(recNum) ;
		roadIceDepth1:long_name = "Road ice depth - sensor 1" ;
		roadIceDepth1:units = "mm" ;
		roadIceDepth1:_FillValue = 3.402823e+38f ;
		roadIceDepth1:missing_value = -9999.f ;
	float roadIceDepth2(recNum) ;
		roadIceDepth2:long_name = "Road ice depth - sensor 2" ;
		roadIceDepth2:units = "mm" ;
		roadIceDepth2:_FillValue = 3.402823e+38f ;
		roadIceDepth2:missing_value = -9999.f ;
	float roadIceDepth3(recNum) ;
		roadIceDepth3:long_name = "Road ice depth - sensor 3" ;
		roadIceDepth3:units = "mm" ;
		roadIceDepth3:_FillValue = 3.402823e+38f ;
		roadIceDepth3:missing_value = -9999.f ;
	float roadIceDepth4(recNum) ;
		roadIceDepth4:long_name = "Road ice depth - sensor 4" ;
		roadIceDepth4:units = "mm" ;
		roadIceDepth4:_FillValue = 3.402823e+38f ;
		roadIceDepth4:missing_value = -9999.f ;
	float roadSnowDepth1(recNum) ;
		roadSnowDepth1:long_name = "Road snow depth - sensor 1" ;
		roadSnowDepth1:units = "cm" ;
		roadSnowDepth1:_FillValue = 3.402823e+38f ;
		roadSnowDepth1:missing_value = -9999.f ;
	float roadSnowDepth2(recNum) ;
		roadSnowDepth2:long_name = "Road snow depth - sensor 2" ;
		roadSnowDepth2:units = "cm" ;
		roadSnowDepth2:_FillValue = 3.402823e+38f ;
		roadSnowDepth2:missing_value = -9999.f ;
	float roadSnowDepth3(recNum) ;
		roadSnowDepth3:long_name = "Road snow depth - sensor 3" ;
		roadSnowDepth3:units = "cm" ;
		roadSnowDepth3:_FillValue = 3.402823e+38f ;
		roadSnowDepth3:missing_value = -9999.f ;
	float roadSnowDepth4(recNum) ;
		roadSnowDepth4:long_name = "Road snow depth - sensor 4" ;
		roadSnowDepth4:units = "cm" ;
		roadSnowDepth4:_FillValue = 3.402823e+38f ;
		roadSnowDepth4:missing_value = -9999.f ;
	float roadLiquidDepth1(recNum) ;
		roadLiquidDepth1:long_name = "Road liquid depth" ;
		roadLiquidDepth1:units = "meter" ;
		roadLiquidDepth1:_FillValue = 3.402823e+38f ;
		roadLiquidDepth1:missing_value = -9999.f ;
	float roadLiquidFreezeTemp1(recNum) ;
		roadLiquidFreezeTemp1:long_name = "Road liquid freezing temp - sensor 1" ;
		roadLiquidFreezeTemp1:units = "kelvin" ;
		roadLiquidFreezeTemp1:_FillValue = 3.402823e+38f ;
		roadLiquidFreezeTemp1:missing_value = -9999.f ;
	float roadLiquidFreezeTemp2(recNum) ;
		roadLiquidFreezeTemp2:long_name = "Road liquid freezing temp - sensor 2" ;
		roadLiquidFreezeTemp2:units = "kelvin" ;
		roadLiquidFreezeTemp2:_FillValue = 3.402823e+38f ;
		roadLiquidFreezeTemp2:missing_value = -9999.f ;
	float roadLiquidFreezeTemp3(recNum) ;
		roadLiquidFreezeTemp3:long_name = "Road liquid freezing temp - sensor 3" ;
		roadLiquidFreezeTemp3:units = "kelvin" ;
		roadLiquidFreezeTemp3:_FillValue = 3.402823e+38f ;
		roadLiquidFreezeTemp3:missing_value = -9999.f ;
	float roadLiquidFreezeTemp4(recNum) ;
		roadLiquidFreezeTemp4:long_name = "Road liquid freezing temp - sensor 4" ;
		roadLiquidFreezeTemp4:units = "kelvin" ;
		roadLiquidFreezeTemp4:_FillValue = 3.402823e+38f ;
		roadLiquidFreezeTemp4:missing_value = -9999.f ;
	float roadLiquidIcePercent1(recNum) ;
		roadLiquidIcePercent1:long_name = "Road liquid ice percent  - sensor 1" ;
		roadLiquidIcePercent1:units = "percent" ;
		roadLiquidIcePercent1:_FillValue = 3.402823e+38f ;
		roadLiquidIcePercent1:missing_value = -9999.f ;
	float roadLiquidIcePercent2(recNum) ;
		roadLiquidIcePercent2:long_name = "Road liquid ice percent  - sensor 2" ;
		roadLiquidIcePercent2:units = "percent" ;
		roadLiquidIcePercent2:_FillValue = 3.402823e+38f ;
		roadLiquidIcePercent2:missing_value = -9999.f ;
	float roadLiquidIcePercent3(recNum) ;
		roadLiquidIcePercent3:long_name = "Road liquid ice percent  - sensor 3" ;
		roadLiquidIcePercent3:units = "percent" ;
		roadLiquidIcePercent3:_FillValue = 3.402823e+38f ;
		roadLiquidIcePercent3:missing_value = -9999.f ;
	float roadLiquidIcePercent4(recNum) ;
		roadLiquidIcePercent4:long_name = "Road liquid ice percent  - sensor 4" ;
		roadLiquidIcePercent4:units = "percent" ;
		roadLiquidIcePercent4:_FillValue = 3.402823e+38f ;
		roadLiquidIcePercent4:missing_value = -9999.f ;

// global attributes:
		:Conventions = "MADIS-like surface observations" ;
		:title = "Built from differnt obs CSV file using csv2madis" ;
}
