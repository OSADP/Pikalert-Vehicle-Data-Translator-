netcdf roads {
dimensions:
	point_num = UNLIMITED ; 
	seg_name_len = 42 ;
	aux_id_len = 8;
	road_type_len = 8 ;
	highway_symbol_len = 8 ;
	num_road_type = 10 ;
	highway_type_len = 1 ;
	rwfs_id_len = 32 ;
variables:
	double latitude(point_num) ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:valid_range = -90., 90. ;
		latitude:units = "degrees_north" ;
	double mid_point_latitude(point_num) ;
		mid_point_latitude:long_name = "latitude of the road segment mid point" ;
		mid_point_latitude:standard_name = "mid point latitude" ;
		mid_point_latitude:valid_range = -90., 90. ;
		mid_point_latitude:units = "degrees_north" ;
	double longitude(point_num) ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:valid_range = -180., 180. ;
		longitude:units = "degrees_east" ;
	double mid_point_longitude(point_num) ;
		mid_point_longitude:long_name = "longitude of the road segment mid point" ;
		mid_point_longitude:standard_name = "mid point longitude" ;
		mid_point_longitude:valid_range = -180., 180. ;
		mid_point_longitude:units = "degrees_east" ;
	float elevation(point_num) ;
		elevation:long_name = "elevation" ;
		elevation:standard_name = "elevation" ;
		elevation:units = "feet" ;
		elevation:_FillValue = -9999.f ;
	char seg_name(point_num, seg_name_len) ;
		seg_name:long_name = "road identifier number for point" ;
		seg_name:standard_name = "road identifier" ;
		seg_name:units = "" ;
	int seg_id(point_num) ;
		seg_id:long_name = "segment identifier for point" ;
		seg_id:standard_name = "segment identifier" ;
	char aux_id(point_num, aux_id_len) ;
		aux_id:long_name = "auxiliary identifier" ;
		aux_id:standard_name = "auxiliary identifier" ;
	int point_type(point_num) ;
		point_type:long_name = "point type" ;
		point_type:flag_values = 0, 1 ;
		point_type:flag_meanings = "road_seg rwis_site" ;
	char rwfs_id(point_num, rwfs_id_len) ;
		rwfs_id:long_name = "corresponding rwfs site id" ;
		rwfs_id:standard_name = "road identifier" ;
	char road_type(point_num, road_type_len) ;
		road_type:long_name = "road type" ;
	short route_class(point_num) ;
		route_class:long_name = "class route" ;
	char highway_type(point_num, highway_type_len) ;
		highway_type:long_name = "highway type" ;
	float speed_mph(point_num) ;
		speed_mph:long_name = "speed miles per hour" ;
		speed_mph:standard_name = "speed_mph" ;
		speed_mph:valid_range = 0., 120. ;
		speed_mph:units = "mi" ;

// global attributes:
		:title = "road segments and rwis sites" ;
		:version = 1. ;
		:Conventions = "CF-1.0" ;
		:description = "" ;
		:observationDimension = "point_num" ;
		:notes = "" ;
}
