netcdf generic_pirep_field_data {

dimensions:
	rec_num = UNLIMITED ; 
	stat_field_name_length = 32;
	num_stat_fields = 40;

variables:

	char stat_field_names(num_stat_fields, stat_field_name_length) ;
	
	double time(rec_num) ;
                time:long_name = "time" ;
                time:units = "seconds since 1970-1-1 00:00" ;
	        
	float latitude(rec_num) ;
		latitude:long_name = "Pirep latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:valid_range = -90., 90. ;
		latitude:units = "degrees_north" ;
		latitude:_FillValue = -99.f ;

	float longitude(rec_num) ;
		longitude:long_name = "Pirep longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:valid_range = -180., 180. ;
		longitude:units = "degrees_east" ;
		longitude:_FillValue = -999.f ;

	int temperature(rec_num) ;
		temperature:long_name = "Temperature" ;
		temperature:units = "degrees C" ;
		temperature:valid_range = -200, 200 ;
		temperature:_FillValue = -999 ;

	byte qpf(rec_num) ;
		qpf:long_name = "Liquid-Equivalent Precipitation Amount" ;
	        qpf:units = "mm tenths" ;

	double mark ;
	        mark:long_name = "bogus" ;


// global attributes:
		:title = "test records" ;
		:version = 1.0 ;
		:Conventions = "CF-1.0" ;
		:description = "" ;
		:observationDimension = "rec_num" ;
		:notes = "" ;

}
